module uart_hw_test (clk,rst_n,txd,rxd);

input clk,rst_n;
input rxd;
output txd;

reg [7:0] tx_data;
reg tx_data_valid;
wire tx_data_ack;
wire txd,rxd;
wire [7:0] rx_data;
wire rx_data_fresh;

reg [7:0] rst_cntr;
reg rst;
always @(posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		rst_cntr <= 0;
		rst <= 1'b1;
	end
	else begin
		if (&rst_cntr) begin
			rst <= 1'b0;
		end
		else begin
			rst <= 1'b1;
			rst_cntr <= rst_cntr + 1'b1;
		end
	end
end

uart u (.clk(clk),
		.rst(rst),
		.tx_data(tx_data),
		.tx_data_valid(tx_data_valid),
		.tx_data_ack(tx_data_ack),
		.txd(txd),
		.rx_data(rx_data),
		.rx_data_fresh(rx_data_fresh),
		.rxd(rxd));

defparam u .CLK_HZ = 100_000_000;
defparam u .BAUD = 115200;

// add one to each RX byte and send it out again
always @(posedge clk) begin
	if (rst) begin
		tx_data <= 1'b0;
		tx_data_valid <= 1'b0;
	end
	else begin
		if (rx_data_fresh) begin
			tx_data <= rx_data + 1'b1;
			tx_data_valid <= 1'b1;
		end	
		else if (tx_data_ack) begin
			tx_data_valid <= 1'b0;
		end
	end
end

endmodule